module spi2axi();
endmodule
